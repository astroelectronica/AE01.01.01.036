.title KiCad schematic
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/C2012CH2A103J125AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C3225X7S1H106M250AB_p.mod"
.include "models/ZXCT1030.spice.txt"
V1 /VIN 0 {VSUPPLY}
XU1 +5V 0 C3225X7S1H106M250AB_p
XU2 +5V 0 C2012X7R2A104K125AA_p
XU4 /CURRENT_FEEDBACK 0 C2012C0G2A102J060AA_p
R5 /CURRENT_FEEDBACK /VOCM 100
V2 +5V 0 5
R6 +5V /TRP 9.76K
R7 /TRP 0 8.66K
R1 /VIN /VOUT 0.47
R2 /VIN /VOUT 0.47
R3 /VOUT /VSN 10K
XU5 /VIN /VSN C2012CH2A103J125AA_p
R4 +5V /ALARM 10K
I1 /VOUT 0 {ILOAD}
XU3 +5V /VSN /VIN 0 /TRP NC_01 /VOCM /ALARM ZXCT1030
.end
